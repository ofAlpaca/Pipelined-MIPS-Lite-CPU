module Shifter(out, B, A);

input [0:31]A, B;
output [0:31]out;

wire [0:31]w1, w2, w3, w4;

TwoToOneMux TTOM10(w1[0], B[31], A[1], A[0]);
TwoToOneMux TTOM11(w1[1], B[31], A[2], A[1]);
TwoToOneMux TTOM12(w1[2], B[31], A[3], A[2]);
TwoToOneMux TTOM13(w1[3], B[31], A[4], A[3]);
TwoToOneMux TTOM14(w1[4], B[31], A[5], A[4]);
TwoToOneMux TTOM15(w1[5], B[31], A[6], A[5]);
TwoToOneMux TTOM16(w1[6], B[31], A[7], A[6]);
TwoToOneMux TTOM17(w1[7], B[31], A[8], A[7]);
TwoToOneMux TTOM18(w1[8], B[31], A[9], A[8]);
TwoToOneMux TTOM19(w1[9], B[31], A[10], A[9]);
TwoToOneMux TTOM110(w1[10], B[31], A[11], A[10]);
TwoToOneMux TTOM111(w1[11], B[31], A[12], A[11]);
TwoToOneMux TTOM112(w1[12], B[31], A[13], A[12]);
TwoToOneMux TTOM113(w1[13], B[31], A[14], A[13]);
TwoToOneMux TTOM114(w1[14], B[31], A[15], A[14]);
TwoToOneMux TTOM115(w1[15], B[31], A[16], A[15]);
TwoToOneMux TTOM116(w1[16], B[31], A[17], A[16]);
TwoToOneMux TTOM117(w1[17], B[31], A[18], A[17]);
TwoToOneMux TTOM118(w1[18], B[31], A[19], A[18]);
TwoToOneMux TTOM119(w1[19], B[31], A[20], A[19]);
TwoToOneMux TTOM120(w1[20], B[31], A[21], A[20]);
TwoToOneMux TTOM121(w1[21], B[31], A[22], A[21]);
TwoToOneMux TTOM122(w1[22], B[31], A[23], A[22]);
TwoToOneMux TTOM123(w1[23], B[31], A[24], A[23]);
TwoToOneMux TTOM124(w1[24], B[31], A[25], A[24]);
TwoToOneMux TTOM125(w1[25], B[31], A[26], A[25]);
TwoToOneMux TTOM126(w1[26], B[31], A[27], A[26]);
TwoToOneMux TTOM127(w1[27], B[31], A[28], A[27]);
TwoToOneMux TTOM128(w1[28], B[31], A[29], A[28]);
TwoToOneMux TTOM129(w1[29], B[31], A[30], A[29]);
TwoToOneMux TTOM130(w1[30], B[31], A[31], A[30]);
TwoToOneMux TTOM131(w1[31], B[31], 1'b0, A[31]);

TwoToOneMux TTOM20(w2[0], B[30], w1[2], w1[0]);
TwoToOneMux TTOM21(w2[1], B[30], w1[3], w1[1]);
TwoToOneMux TTOM22(w2[2], B[30], w1[4], w1[2]);
TwoToOneMux TTOM23(w2[3], B[30], w1[5], w1[3]);
TwoToOneMux TTOM24(w2[4], B[30], w1[6], w1[4]);
TwoToOneMux TTOM25(w2[5], B[30], w1[7], w1[5]);
TwoToOneMux TTOM26(w2[6], B[30], w1[8], w1[6]);
TwoToOneMux TTOM27(w2[7], B[30], w1[9], w1[7]);
TwoToOneMux TTOM28(w2[8], B[30], w1[10], w1[8]);
TwoToOneMux TTOM29(w2[9], B[30], w1[11], w1[9]);
TwoToOneMux TTOM210(w2[10], B[30], w1[12], w1[10]);
TwoToOneMux TTOM211(w2[11], B[30], w1[13], w1[11]);
TwoToOneMux TTOM212(w2[12], B[30], w1[14], w1[12]);
TwoToOneMux TTOM213(w2[13], B[30], w1[15], w1[13]);
TwoToOneMux TTOM214(w2[14], B[30], w1[16], w1[14]);
TwoToOneMux TTOM215(w2[15], B[30], w1[17], w1[15]);
TwoToOneMux TTOM216(w2[16], B[30], w1[18], w1[16]);
TwoToOneMux TTOM217(w2[17], B[30], w1[19], w1[17]);
TwoToOneMux TTOM218(w2[18], B[30], w1[20], w1[18]);
TwoToOneMux TTOM219(w2[19], B[30], w1[21], w1[19]);
TwoToOneMux TTOM220(w2[20], B[30], w1[22], w1[20]);
TwoToOneMux TTOM221(w2[21], B[30], w1[23], w1[21]);
TwoToOneMux TTOM222(w2[22], B[30], w1[24], w1[22]);
TwoToOneMux TTOM223(w2[23], B[30], w1[25], w1[23]);
TwoToOneMux TTOM224(w2[24], B[30], w1[26], w1[24]);
TwoToOneMux TTOM225(w2[25], B[30], w1[27], w1[25]);
TwoToOneMux TTOM226(w2[26], B[30], w1[28], w1[26]);
TwoToOneMux TTOM227(w2[27], B[30], w1[29], w1[27]);
TwoToOneMux TTOM228(w2[28], B[30], w1[30], w1[28]);
TwoToOneMux TTOM229(w2[29], B[30], w1[31], w1[29]);
TwoToOneMux TTOM230(w2[30], B[30], 1'b0, w1[30]);
TwoToOneMux TTOM231(w2[31], B[30], 1'b0, w1[31]);

TwoToOneMux TTOM30(w3[0], B[29], w2[4], w2[0]);
TwoToOneMux TTOM31(w3[1], B[29], w2[5], w2[1]);
TwoToOneMux TTOM32(w3[2], B[29], w2[6], w2[2]);
TwoToOneMux TTOM33(w3[3], B[29], w2[7], w2[3]);
TwoToOneMux TTOM34(w3[4], B[29], w2[8], w2[4]);
TwoToOneMux TTOM35(w3[5], B[29], w2[9], w2[5]);
TwoToOneMux TTOM36(w3[6], B[29], w2[10], w2[6]);
TwoToOneMux TTOM37(w3[7], B[29], w2[11], w2[7]);
TwoToOneMux TTOM38(w3[8], B[29], w2[12], w2[8]);
TwoToOneMux TTOM39(w3[9], B[29], w2[13], w2[9]);
TwoToOneMux TTOM310(w3[10], B[29], w2[14], w2[10]);
TwoToOneMux TTOM311(w3[11], B[29], w2[15], w2[11]);
TwoToOneMux TTOM312(w3[12], B[29], w2[16], w2[12]);
TwoToOneMux TTOM313(w3[13], B[29], w2[17], w2[13]);
TwoToOneMux TTOM314(w3[14], B[29], w2[18], w2[14]);
TwoToOneMux TTOM315(w3[15], B[29], w2[19], w2[15]);
TwoToOneMux TTOM316(w3[16], B[29], w2[20], w2[16]);
TwoToOneMux TTOM317(w3[17], B[29], w2[21], w2[17]);
TwoToOneMux TTOM318(w3[18], B[29], w2[22], w2[18]);
TwoToOneMux TTOM319(w3[19], B[29], w2[23], w2[19]);
TwoToOneMux TTOM320(w3[20], B[29], w2[24], w2[20]);
TwoToOneMux TTOM321(w3[21], B[29], w2[25], w2[21]);
TwoToOneMux TTOM322(w3[22], B[29], w2[26], w2[22]);
TwoToOneMux TTOM323(w3[23], B[29], w2[27], w2[23]);
TwoToOneMux TTOM324(w3[24], B[29], w2[28], w2[24]);
TwoToOneMux TTOM325(w3[25], B[29], w2[29], w2[25]);
TwoToOneMux TTOM326(w3[26], B[29], w2[30], w2[26]);
TwoToOneMux TTOM327(w3[27], B[29], w2[31], w2[27]);
TwoToOneMux TTOM328(w3[28], B[29], 1'b0, w2[28]);
TwoToOneMux TTOM329(w3[29], B[29], 1'b0, w2[29]);
TwoToOneMux TTOM330(w3[30], B[29], 1'b0, w2[30]);
TwoToOneMux TTOM331(w3[31], B[29], 1'b0, w2[31]);

TwoToOneMux TTOM40(w4[0], B[28], w3[8], w3[0]);
TwoToOneMux TTOM41(w4[1], B[28], w3[9], w3[1]);
TwoToOneMux TTOM42(w4[2], B[28], w3[10], w3[2]);
TwoToOneMux TTOM43(w4[3], B[28], w3[11], w3[3]);
TwoToOneMux TTOM44(w4[4], B[28], w3[12], w3[4]);
TwoToOneMux TTOM45(w4[5], B[28], w3[13], w3[5]);
TwoToOneMux TTOM46(w4[6], B[28], w3[14], w3[6]);
TwoToOneMux TTOM47(w4[7], B[28], w3[15], w3[7]);
TwoToOneMux TTOM48(w4[8], B[28], w3[16], w3[8]);
TwoToOneMux TTOM49(w4[9], B[28], w3[17], w3[9]);
TwoToOneMux TTOM410(w4[10], B[28], w3[18], w3[10]);
TwoToOneMux TTOM411(w4[11], B[28], w3[19], w3[11]);
TwoToOneMux TTOM412(w4[12], B[28], w3[20], w3[12]);
TwoToOneMux TTOM413(w4[13], B[28], w3[21], w3[13]);
TwoToOneMux TTOM414(w4[14], B[28], w3[22], w3[14]);
TwoToOneMux TTOM415(w4[15], B[28], w3[23], w3[15]);
TwoToOneMux TTOM416(w4[16], B[28], w3[24], w3[16]);
TwoToOneMux TTOM417(w4[17], B[28], w3[25], w3[17]);
TwoToOneMux TTOM418(w4[18], B[28], w3[26], w3[18]);
TwoToOneMux TTOM419(w4[19], B[28], w3[27], w3[19]);
TwoToOneMux TTOM420(w4[20], B[28], w3[28], w3[20]);
TwoToOneMux TTOM421(w4[21], B[28], w3[29], w3[21]);
TwoToOneMux TTOM422(w4[22], B[28], w3[30], w3[22]);
TwoToOneMux TTOM423(w4[23], B[28], w3[31], w3[23]);
TwoToOneMux TTOM424(w4[24], B[28], 1'b0, w3[24]);
TwoToOneMux TTOM425(w4[25], B[28], 1'b0, w3[25]);
TwoToOneMux TTOM426(w4[26], B[28], 1'b0, w3[26]);
TwoToOneMux TTOM427(w4[27], B[28], 1'b0, w3[27]);
TwoToOneMux TTOM428(w4[28], B[28], 1'b0, w3[28]);
TwoToOneMux TTOM429(w4[29], B[28], 1'b0, w3[29]);
TwoToOneMux TTOM430(w4[30], B[28], 1'b0, w3[30]);
TwoToOneMux TTOM431(w4[31], B[28], 1'b0, w3[31]);

TwoToOneMux TTOM50(out[0], B[27], w4[16], w4[0]);
TwoToOneMux TTOM51(out[1], B[27], w4[17], w4[1]);
TwoToOneMux TTOM52(out[2], B[27], w4[18], w4[2]);
TwoToOneMux TTOM53(out[3], B[27], w4[19], w4[3]);
TwoToOneMux TTOM54(out[4], B[27], w4[20], w4[4]);
TwoToOneMux TTOM55(out[5], B[27], w4[21], w4[5]);
TwoToOneMux TTOM56(out[6], B[27], w4[22], w4[6]);
TwoToOneMux TTOM57(out[7], B[27], w4[23], w4[7]);
TwoToOneMux TTOM58(out[8], B[27], w4[24], w4[8]);
TwoToOneMux TTOM59(out[9], B[27], w4[25], w4[9]);
TwoToOneMux TTOM510(out[10], B[27], w4[26], w4[10]);
TwoToOneMux TTOM511(out[11], B[27], w4[27], w4[11]);
TwoToOneMux TTOM512(out[12], B[27], w4[28], w4[12]);
TwoToOneMux TTOM513(out[13], B[27], w4[29], w4[13]);
TwoToOneMux TTOM514(out[14], B[27], w4[30], w4[14]);
TwoToOneMux TTOM515(out[15], B[27], w4[31], w4[15]);
TwoToOneMux TTOM516(out[16], B[27], 1'b0, w4[16]);
TwoToOneMux TTOM517(out[17], B[27], 1'b0, w4[17]);
TwoToOneMux TTOM518(out[18], B[27], 1'b0, w4[18]);
TwoToOneMux TTOM519(out[19], B[27], 1'b0, w4[19]);
TwoToOneMux TTOM520(out[20], B[27], 1'b0, w4[20]);
TwoToOneMux TTOM521(out[21], B[27], 1'b0, w4[21]);
TwoToOneMux TTOM522(out[22], B[27], 1'b0, w4[22]);
TwoToOneMux TTOM523(out[23], B[27], 1'b0, w4[23]);
TwoToOneMux TTOM524(out[24], B[27], 1'b0, w4[24]);
TwoToOneMux TTOM525(out[25], B[27], 1'b0, w4[25]);
TwoToOneMux TTOM526(out[26], B[27], 1'b0, w4[26]);
TwoToOneMux TTOM527(out[27], B[27], 1'b0, w4[27]);
TwoToOneMux TTOM528(out[28], B[27], 1'b0, w4[28]);
TwoToOneMux TTOM529(out[29], B[27], 1'b0, w4[29]);
TwoToOneMux TTOM530(out[30], B[27], 1'b0, w4[30]);
TwoToOneMux TTOM531(out[31], B[27], 1'b0, w4[31]);

endmodule
